`define INWVAL 12
`define RVAL 9
`define CVAL 8
`define MAXKVAL 5
`define TVPR 0.65
`define TRPR 0.7
