`define INWVAL 24
`define RVAL 16
`define CVAL 17
`define MAXKVAL 9
`define TVPR 1.0
`define TRPR 1.0
