`define INWVAL 18
`define RVAL 9
`define CVAL 8
`define MAXKVAL 5
`define TVPR 1.0
`define TRPR 1.0
