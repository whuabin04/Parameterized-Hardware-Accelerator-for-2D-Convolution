`define INWVAL 12
`define OUTWVAL 24
`define PIPELINEDVAL 1
